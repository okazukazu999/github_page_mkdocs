name: Deploy mkdocs

on:
  pull_request:
    # PRのcloseをトリガーとしてjobを実行する
    branches:
      - master
    types:
      - closed

jobs:
  deploy:
    runs-on: ubuntu-18.04
    steps:

      - run: echo "Hello, World!"



      - name: checkout branch 
        uses: actions/checkout@v2
        with:
          fetch-depth: 0

      - name: configure git info
        run: |
          git config --global user.name "github-actions-for-deploy"
          git config --global user.email deploy-actions@github.com
      - name: check git status/branch
        run: |
          git status
          git branch
      # mkdocsを利用するためのpython環境のセットアップ
      - name: setup python env
        uses: actions/setup-python@v1
        with:
          python-version: '3.8'

      - name: install dependencies
        run: |
          # python -m pip install --upgrade pip
          pip install -r requirements.txt
      # ドキュメントの作成
      - name: mkdocs build
        run: |
           mkdocs build --verbose --clean --strict
      # ドキュメントのデプロイ
      - name: mkdocs deploy
        uses: peaceiris/actions-gh-pages@v3
        with:
           github_token: ${{ secrets.PERSONAL_TOKEN }}
           publish_dir: site
